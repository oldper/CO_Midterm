`include "mux_2to1.v"
module Shifter( dataA, shamt, Signal, dataOut);
input reset ;
input [31:0] dataA ;
input [5:0] shamt;
input [4:0] Signal ;
output [31:0] dataOut ;

parameter SRL = 6'b000010;


wire [31:0] wire1;
wire [31:0] wire2;
wire [31:0] wire3;
wire [31:0] wire4;
wire [31:0] wire5;

mux_2to1 m000( wire1[0], dataA[0], dataA[1], shamt[0] );
mux_2to1 m001( wire1[1], dataA[1], dataA[2], shamt[0] );
mux_2to1 m002( wire1[2], dataA[2], dataA[3], shamt[0] );
mux_2to1 m003( wire1[3], dataA[3], dataA[4], shamt[0] );
mux_2to1 m004( wire1[4], dataA[4], dataA[5], shamt[0] );
mux_2to1 m005( wire1[5], dataA[5], dataA[6], shamt[0] );
mux_2to1 m006( wire1[6], dataA[6], dataA[7], shamt[0] );
mux_2to1 m007( wire1[7], dataA[7], dataA[8], shamt[0] );
mux_2to1 m008( wire1[8], dataA[8], dataA[9], shamt[0] );
mux_2to1 m009( wire1[9], dataA[9], dataA[10], shamt[0] );
mux_2to1 m010( wire1[10], dataA[10], dataA[11], shamt[0] );
mux_2to1 m011( wire1[11], dataA[11], dataA[12], shamt[0] );
mux_2to1 m012( wire1[12], dataA[12], dataA[13], shamt[0] );
mux_2to1 m013( wire1[13], dataA[13], dataA[14], shamt[0] );
mux_2to1 m014( wire1[14], dataA[14], dataA[15], shamt[0] );
mux_2to1 m015( wire1[15], dataA[15], dataA[16], shamt[0] );
mux_2to1 m016( wire1[16], dataA[16], dataA[17], shamt[0] );
mux_2to1 m017( wire1[17], dataA[17], dataA[18], shamt[0] );
mux_2to1 m018( wire1[18], dataA[18], dataA[19], shamt[0] );
mux_2to1 m019( wire1[19], dataA[19], dataA[20], shamt[0] );
mux_2to1 m020( wire1[20], dataA[20], dataA[21], shamt[0] );
mux_2to1 m021( wire1[21], dataA[21], dataA[22], shamt[0] );
mux_2to1 m022( wire1[22], dataA[22], dataA[23], shamt[0] );
mux_2to1 m023( wire1[23], dataA[23], dataA[24], shamt[0] );
mux_2to1 m024( wire1[24], dataA[24], dataA[25], shamt[0] );
mux_2to1 m025( wire1[25], dataA[25], dataA[26], shamt[0] );
mux_2to1 m026( wire1[26], dataA[26], dataA[27], shamt[0] );
mux_2to1 m027( wire1[27], dataA[27], dataA[28], shamt[0] );
mux_2to1 m028( wire1[28], dataA[28], dataA[29], shamt[0] );
mux_2to1 m029( wire1[29], dataA[29], dataA[30], shamt[0] );
mux_2to1 m030( wire1[30], dataA[30], dataA[31], shamt[0] );
mux_2to1 m031( wire1[31], dataA[31], 1'b0, shamt[0] );

mux_2to1 m100( wire2[0], wire1[0], wire1[2], shamt[1] );
mux_2to1 m101( wire2[1], wire1[1], wire1[3], shamt[1] );
mux_2to1 m102( wire2[2], wire1[2], wire1[4], shamt[1] );
mux_2to1 m103( wire2[3], wire1[3], wire1[5], shamt[1] );
mux_2to1 m104( wire2[4], wire1[4], wire1[6], shamt[1] );
mux_2to1 m105( wire2[5], wire1[5], wire1[7], shamt[1] );
mux_2to1 m106( wire2[6], wire1[6], wire1[8], shamt[1] );
mux_2to1 m107( wire2[7], wire1[7], wire1[9], shamt[1] );
mux_2to1 m108( wire2[8], wire1[8], wire1[10], shamt[1] );
mux_2to1 m109( wire2[9], wire1[9], wire1[11], shamt[1] );
mux_2to1 m110( wire2[10], wire1[10], wire1[12], shamt[1] );
mux_2to1 m111( wire2[11], wire1[11], wire1[13], shamt[1] );
mux_2to1 m112( wire2[12], wire1[12], wire1[14], shamt[1] );
mux_2to1 m113( wire2[13], wire1[13], wire1[15], shamt[1] );
mux_2to1 m114( wire2[14], wire1[14], wire1[16], shamt[1] );
mux_2to1 m115( wire2[15], wire1[15], wire1[17], shamt[1] );
mux_2to1 m116( wire2[16], wire1[16], wire1[18], shamt[1] );
mux_2to1 m117( wire2[17], wire1[17], wire1[19], shamt[1] );
mux_2to1 m118( wire2[18], wire1[18], wire1[20], shamt[1] );
mux_2to1 m119( wire2[19], wire1[19], wire1[21], shamt[1] );
mux_2to1 m120( wire2[20], wire1[20], wire1[22], shamt[1] );
mux_2to1 m121( wire2[21], wire1[21], wire1[23], shamt[1] );
mux_2to1 m122( wire2[22], wire1[22], wire1[24], shamt[1] );
mux_2to1 m123( wire2[23], wire1[23], wire1[25], shamt[1] );
mux_2to1 m124( wire2[24], wire1[24], wire1[26], shamt[1] );
mux_2to1 m125( wire2[25], wire1[25], wire1[27], shamt[1] );
mux_2to1 m126( wire2[26], wire1[26], wire1[28], shamt[1] );
mux_2to1 m127( wire2[27], wire1[27], wire1[29], shamt[1] );
mux_2to1 m128( wire2[28], wire1[28], wire1[30], shamt[1] );
mux_2to1 m129( wire2[29], wire1[29], wire1[31], shamt[1] );
mux_2to1 m130( wire2[30], wire1[30], 1'b0, shamt[1] );
mux_2to1 m131( wire2[31], wire1[31], 1'b0, shamt[1] );


mux_2to1 m200( wire3[0], wire2[0], wire2[4], shamt[2] );
mux_2to1 m201( wire3[1], wire2[1], wire2[5], shamt[2] );
mux_2to1 m202( wire3[2], wire2[2], wire2[6], shamt[2] );
mux_2to1 m203( wire3[3], wire2[3], wire2[7], shamt[2] );
mux_2to1 m204( wire3[4], wire2[4], wire2[8], shamt[2] );
mux_2to1 m205( wire3[5], wire2[5], wire2[9], shamt[2] );
mux_2to1 m206( wire3[6], wire2[6], wire2[10], shamt[2] );
mux_2to1 m207( wire3[7], wire2[7], wire2[11], shamt[2] );
mux_2to1 m208( wire3[8], wire2[8], wire2[12], shamt[2] );
mux_2to1 m209( wire3[9], wire2[9], wire2[13], shamt[2] );
mux_2to1 m210( wire3[10], wire2[10], wire2[14], shamt[2] );
mux_2to1 m211( wire3[11], wire2[11], wire2[15], shamt[2] );
mux_2to1 m212( wire3[12], wire2[12], wire2[16], shamt[2] );
mux_2to1 m213( wire3[13], wire2[13], wire2[17], shamt[2] );
mux_2to1 m214( wire3[14], wire2[14], wire2[18], shamt[2] );
mux_2to1 m215( wire3[15], wire2[15], wire2[19], shamt[2] );
mux_2to1 m216( wire3[16], wire2[16], wire2[20], shamt[2] );
mux_2to1 m217( wire3[17], wire2[17], wire2[21], shamt[2] );
mux_2to1 m218( wire3[18], wire2[18], wire2[22], shamt[2] );
mux_2to1 m219( wire3[19], wire2[19], wire2[23], shamt[2] );
mux_2to1 m220( wire3[20], wire2[20], wire2[24], shamt[2] );
mux_2to1 m221( wire3[21], wire2[21], wire2[25], shamt[2] );
mux_2to1 m222( wire3[22], wire2[22], wire2[26], shamt[2] );
mux_2to1 m223( wire3[23], wire2[23], wire2[27], shamt[2] );
mux_2to1 m224( wire3[24], wire2[24], wire2[28], shamt[2] );
mux_2to1 m225( wire3[25], wire2[25], wire2[29], shamt[2] );
mux_2to1 m226( wire3[26], wire2[26], wire2[30], shamt[2] );
mux_2to1 m227( wire3[27], wire2[27], wire2[31], shamt[2] );
mux_2to1 m228( wire3[28], wire2[28], 1'b0, shamt[2] );
mux_2to1 m229( wire3[29], wire2[29], 1'b0, shamt[2] );
mux_2to1 m230( wire3[30], wire2[30], 1'b0, shamt[2] );
mux_2to1 m231( wire3[31], wire2[31], 1'b0, shamt[2] );

mux_2to1 m300( wire4[0], wire3[0], wire3[8], shamt[3] );
mux_2to1 m301( wire4[1], wire3[1], wire3[9], shamt[3] );
mux_2to1 m302( wire4[2], wire3[2], wire3[10], shamt[3] );
mux_2to1 m303( wire4[3], wire3[3], wire3[11], shamt[3] );
mux_2to1 m304( wire4[4], wire3[4], wire3[12], shamt[3] );
mux_2to1 m305( wire4[5], wire3[5], wire3[13], shamt[3] );
mux_2to1 m306( wire4[6], wire3[6], wire3[14], shamt[3] );
mux_2to1 m307( wire4[7], wire3[7], wire3[15], shamt[3] );
mux_2to1 m308( wire4[8], wire3[8], wire3[16], shamt[3] );
mux_2to1 m309( wire4[9], wire3[9], wire3[17], shamt[3] );
mux_2to1 m310( wire4[10], wire3[10], wire3[18], shamt[3] );
mux_2to1 m311( wire4[11], wire3[11], wire3[19], shamt[3] );
mux_2to1 m312( wire4[12], wire3[12], wire3[20], shamt[3] );
mux_2to1 m313( wire4[13], wire3[13], wire3[21], shamt[3] );
mux_2to1 m314( wire4[14], wire3[14], wire3[22], shamt[3] );
mux_2to1 m315( wire4[15], wire3[15], wire3[23], shamt[3] );
mux_2to1 m316( wire4[16], wire3[16], wire3[24], shamt[3] );
mux_2to1 m317( wire4[17], wire3[17], wire3[25], shamt[3] );
mux_2to1 m318( wire4[18], wire3[18], wire3[26], shamt[3] );
mux_2to1 m319( wire4[19], wire3[19], wire3[27], shamt[3] );
mux_2to1 m320( wire4[20], wire3[20], wire3[28], shamt[3] );
mux_2to1 m321( wire4[21], wire3[21], wire3[29], shamt[3] );
mux_2to1 m322( wire4[22], wire3[22], wire3[30], shamt[3] );
mux_2to1 m323( wire4[23], wire3[23], wire3[31], shamt[3] );
mux_2to1 m324( wire4[24], wire3[24], 1'b0, shamt[3] );
mux_2to1 m325( wire4[25], wire3[25], 1'b0, shamt[3] );
mux_2to1 m326( wire4[26], wire3[26], 1'b0, shamt[3] );
mux_2to1 m327( wire4[27], wire3[27], 1'b0, shamt[3] );
mux_2to1 m328( wire4[28], wire3[28], 1'b0, shamt[3] );
mux_2to1 m329( wire4[29], wire3[29], 1'b0, shamt[3] );
mux_2to1 m330( wire4[30], wire3[30], 1'b0, shamt[3] );
mux_2to1 m331( wire4[31], wire3[31], 1'b0, shamt[3] );

mux_2to1 m400( dataOut[0], wire4[0], wire4[16], shamt[4] );
mux_2to1 m401( dataOut[1], wire4[1], wire4[17], shamt[4] );
mux_2to1 m402( dataOut[2], wire4[2], wire4[18], shamt[4] );
mux_2to1 m403( dataOut[3], wire4[3], wire4[19], shamt[4] );
mux_2to1 m404( dataOut[4], wire4[4], wire4[20], shamt[4] );
mux_2to1 m405( dataOut[5], wire4[5], wire4[21], shamt[4] );
mux_2to1 m406( dataOut[6], wire4[6], wire4[22], shamt[4] );
mux_2to1 m407( dataOut[7], wire4[7], wire4[23], shamt[4] );
mux_2to1 m408( dataOut[8], wire4[8], wire4[24], shamt[4] );
mux_2to1 m409( dataOut[9], wire4[9], wire4[25], shamt[4] );
mux_2to1 m410( dataOut[10], wire4[10], wire4[26], shamt[4] );
mux_2to1 m411( dataOut[11], wire4[11], wire4[27], shamt[4] );
mux_2to1 m412( dataOut[12], wire4[12], wire4[28], shamt[4] );
mux_2to1 m413( dataOut[13], wire4[13], wire4[29], shamt[4] );
mux_2to1 m414( dataOut[14], wire4[14], wire4[30], shamt[4] );
mux_2to1 m415( dataOut[15], wire4[15], wire4[31], shamt[4] );
mux_2to1 m416( dataOut[16], wire4[16], 1'b0, shamt[4] );
mux_2to1 m417( dataOut[17], wire4[17], 1'b0, shamt[4] );
mux_2to1 m418( dataOut[18], wire4[18], 1'b0, shamt[4] );
mux_2to1 m419( dataOut[19], wire4[19], 1'b0, shamt[4] );
mux_2to1 m420( dataOut[20], wire4[20], 1'b0, shamt[4] );
mux_2to1 m421( dataOut[21], wire4[21], 1'b0, shamt[4] );
mux_2to1 m422( dataOut[22], wire4[22], 1'b0, shamt[4] );
mux_2to1 m423( dataOut[23], wire4[23], 1'b0, shamt[4] );
mux_2to1 m424( dataOut[24], wire4[24], 1'b0, shamt[4] );
mux_2to1 m425( dataOut[25], wire4[25], 1'b0, shamt[4] );
mux_2to1 m426( dataOut[26], wire4[26], 1'b0, shamt[4] );
mux_2to1 m427( dataOut[27], wire4[27], 1'b0, shamt[4] );
mux_2to1 m428( dataOut[28], wire4[28], 1'b0, shamt[4] );
mux_2to1 m429( dataOut[29], wire4[29], 1'b0, shamt[4] );
mux_2to1 m430( dataOut[30], wire4[30], 1'b0, shamt[4] );
mux_2to1 m431( dataOut[31], wire4[31], 1'b0, shamt[4] );

endmodule